module mux2(
    a,
    b,
    s,
    f
);

assign f = (s)?b:a;endmoudle
